----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 31.01.2024 10:44:20
-- Design Name: 
-- Module Name: float_to_int - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
entity left_shift is
    Port (  input: in std_logic_vector(7 downto 0);
            output: out std_logic_vector(7 downto 0);
            samt: in std_logic_vector(3 downto 0));

end left_shift;

architecture Behavioral of left_shift is

begin


end Behavioral;

entity float_to_int is
--  Port ( );
end float_to_int;

architecture Behavioral of float_to_int is

begin


end Behavioral;
